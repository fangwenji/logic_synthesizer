module TestCase2 (input c, input b, output t);
  input c;
  input b;
  output t;
  assign t = b;
endmodule
